/**
 * @file udp_output_header_bfm.sv
 * 
 * @author Mani Magnusson
 * @date   2024
 * 
 * @brief UDP Header (logic to PHY) bus functional model
 */

`timescale 1ns / 1ps
`default_nettype none



`default_nettype wire