/**
 * @file axi-lite_if.sv
 *
 * @author Mani Magnusson
 * @date   2023
 *
 * @brief AXI4-Lite Interface Definition, uses a 32 bit bus
 */

 /*
  * TODO:
  *  - Add this shi
  */

  `default_nettype none

  interface AXIS_IF # ();
  // Signals




  `default_nettype wire