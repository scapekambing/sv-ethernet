/**
 * @file udp_tx_header_bfm.sv
 * 
 * @author Mani Magnusson
 * @date   2024
 * 
 * @brief UDP TX Header (logic to PHY) bus functional model
 */

`timescale 1ns / 1ps
`default_nettype none

package udp_tx_header_bfm;
class UDP_TX_HEADER_SLAVE_BFM # (
    // Parameters
);
    // Do stuff
endclass

class UDP_TX_HEADER_MASTER_BFM # (
    // Parameters
);
    // Do stuff
endclass
endpackage

`default_nettype wire