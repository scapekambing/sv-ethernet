/**
 * @file udp_input_header_bfm.sv
 * 
 * @author Mani Magnusson
 * @date   2024
 * 
 * @brief UDP Header (PHY to logic) bus functional model
 */

`timescale 1ns / 1ps
`default_nettype none



`default_nettype wire