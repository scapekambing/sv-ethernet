/**
 * @file eth_top.sv
 *
 * @author Mani Magnusson
 * @date   2024
 *
 * @brief Top module of Ethernet stack
 */

 `default_nettype none

 module eth_top # (
    // Parameters
 ) (
    // Signals
 );
    // Logic
 endmodule

 `default_nettype wire